module Task7_Cordic_Pipline_top(